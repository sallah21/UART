`timescale 1ns / 100ps
module RX_tb;



endmodule